netcdf mom6_vgrid {
dimensions:
	Layer = 41 ;
	interfaces = 42 ;
variables:
	double dz(Layer) ;
		dz:units = "m" ;
		dz:long_name = "z* coordinate level thickness" ;
	double sigma2(interfaces) ;
		sigma2:units = "kg/m3" ;
		sigma2:long_name = "Interface target potential density references to 2000 dbars" ;
	double Layer(Layer) ;
		Layer:units = "kg/m3" ;
		Layer:long_name = "Layer target potential density references to 2000 dbars" ;
data:

 dz = 1, 1.8, 3.24, 4.68, 4.93, 5.81, 6.87, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 
    8, 8, 8, 8, 8, 10, 16.4, 35.92, 42.38, 50.02, 59.02, 69.64, 82.18, 96.97, 
    114.43, 135.02, 159.33, 188.01, 221.84, 261.78, 400, 600, 600 ;

 sigma2 = 1007, 1011.5, 1014.5, 1018, 1020.5, 1021.5, 1022.5, 1023.5, 1024.5, 
    1025.5, 1026.5, 1027.5, 1028.5, 1029.45, 1030.275, 1031, 1031.65, 
    1032.25, 1032.85, 1033.45, 1034.025, 1034.55, 1035, 1035.35, 1035.65, 
    1035.92, 1036.12, 1036.29, 1036.45, 1036.57, 1036.66, 1036.735, 1036.8, 
    1036.86, 1036.93, 1036.995, 1037.04, 1037.08, 1037.135, 1037.235, 
    1037.36, 1037.54 ;

 Layer = 1010, 1013, 1016, 1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 
    1028, 1029, 1029.9, 1030.65, 1031.35, 1031.95, 1032.55, 1033.15, 1033.75, 
    1034.3, 1034.8, 1035.2, 1035.5, 1035.8, 1036.04, 1036.2, 1036.38, 
    1036.52, 1036.62, 1036.7, 1036.77, 1036.83, 1036.89, 1036.97, 1037.02, 
    1037.06, 1037.1, 1037.17, 1037.3, 1037.42 ;
}
